module plic (
    output bit irq_ext = 1'b0
);
    
endmodule