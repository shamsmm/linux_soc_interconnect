module plic (
    
);
    
endmodule